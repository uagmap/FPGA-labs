-- add necessary libraries and packages
library ieee;
library ieee_proposed;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee_proposed.fixed_float_types.all;
use ieee_proposed.fixed_pkg.all;

entity filter_fsm is
		generic(
					m : natural := 4; -- Qm.n
					n : natural := 12); -- Qm.n
		port( 
			rst           : in  std_logic;
			clk           : in  std_logic;
			enhance       : in  std_logic;
         left_right    : in  std_logic;
         codec_idle    : in  std_logic;
         left_in       : in  std_logic_vector(15 downto 0);
         right_in      : in  std_logic_vector(15 downto 0);
         codec_start   : out std_logic;
         reg_addr      : out std_logic_vector(6 downto 0);
         reg_data      : out std_logic_vector(8 downto 0);
         left_out      : out std_logic_vector(15 downto 0);
         right_out     : out std_logic_vector(15 downto 0)
				);
end filter_fsm;

architecture behavioral of filter_fsm is
    type TState is (idle, config0, wait0, wait1, config1, filter0);
    signal state : TState;
    signal left_right_1 : std_logic;
    constant ROM_SIZE : natural := 9;

    type memory is array (NATURAL range 0 to ROM_SIZE - 1) of std_logic_vector(15 downto 0);
    constant config_rom : memory := (
												"0001111000000000", -- Reset reg.
												"0000111000000010", -- Digital Audio Interface Format reg.
												"0000101000010001", -- Digital Audio Path Control reg.
												"0001000000100011", -- Sampling Control reg. (44.1 kHz, USB mode)
												"0001001000000001", -- Active reg.
												"0000100000010000", -- Analogue Audio Path Control reg.
												"0000110000000000", -- Power Down Control reg.
												"0000000000011000", -- Left Line In reg.
												"0000001000011000"); -- Right Line In reg.

    TYPE delay_line IS ARRAY(0 TO 2) OF SFIXED(m - 1 downto -n);
    TYPE coeff_line IS ARRAY(0 TO 2) OF SFIXED(m - 1 downto -n);

--    constant a : coeff_line := (
--        TO_SFIXED(1.000, m - 1, -n), -- denominator coeff.
--        TO_SFIXED(-1.601092394183619, m - 1, -n),
--        TO_SFIXED(0.668368994611848, m - 1, -n)
--    );
--
--    constant b : coeff_line := (
--        TO_SFIXED(3.269461388795467, m - 1, -n), -- numerator coeff.
--        TO_SFIXED(-6.538922777590933, m - 1, -n),
--        TO_SFIXED(3.269461388795467, m - 1, -n)
--    );


--LOW PASS BELOW
		constant a : coeff_line := (
			  TO_SFIXED(1.000, m - 1, -n), -- denominator coeff.
			  TO_SFIXED(-1.799096409484668, m - 1, -n),
			  TO_SFIXED(0.817512403384758, m - 1, -n)
		 );

		 constant b : coeff_line := (
			  TO_SFIXED(0.018415993900090, m - 1, -n), -- numerator coeff.
			  TO_SFIXED(0.036831987800180, m - 1, -n),
			  TO_SFIXED(0.018415993900090, m - 1, -n)
		 );

    signal z_left, z_right : SFIXED(m downto -n); -- m+n+1 bits to provide space for + oper.
    signal left_out_int : std_logic_vector(m + n downto 0); -- m+n+1 bits to provide space for + oper.
    signal right_out_int : std_logic_vector(m + n downto 0); -- m+n+1 bits to provide space for + oper.

BEGIN
    PROCESS(clk, rst)
        variable rom_ptr : natural := 0;
        variable ram_ptr : natural := 0;
        variable data_reg : std_logic_vector(15 downto 0);
		  
        variable x_left, x_right : delay_line; -- inputs in SFIXED format
        variable y_left, y_right : delay_line; -- output of the trebble filters
        variable acc_left : SFIXED(2 * m - 1 + 4 downto -(2 * n)); -- larger dynamic range for + and * oper.
        variable acc_right : SFIXED(2 * m - 1 + 4 downto -(2 * n)); -- larger dynamic range for + and * oper.
    BEGIN
        IF (rst = '0') THEN
            -- reset signals and variables
				state <= idle;
				left_right_1 <= '0';
				state <= idle;
				rom_ptr := 0;
				ram_ptr := 0;
				codec_start <= '0';
				left_out <= (others => '0');--reset outputs
				right_out <= (others => '0');
				
        ELSIF (clk'EVENT AND clk = '1') THEN
            CASE State IS
               WHEN idle =>
							state <= config0;
					 
               WHEN config0 =>  -- read codec config. info from ROM
                    data_reg := config_rom(rom_ptr); 
                    reg_addr <= data_reg(15 downto 9); -- first seven bits are address
                    reg_data <= data_reg(8 downto 0);
                    codec_start <= '1';
                    state <= wait0;

                WHEN wait0 =>  -- wait until i2c_codec starts transmission
                    IF (codec_idle = '1') THEN
                        state <= wait0;
                    ELSE
                        state <= wait1;
                    END IF;

                WHEN wait1 =>  -- wait for i2c_codec to finish transmission
                    IF (codec_idle = '0') THEN
                        state <= wait1;
                        codec_start <= '0'; --clear start signal
                    ELSE
                        state <= config1;
                    END IF;

                WHEN config1 =>  -- check if ROM has been fully read
                    rom_ptr := rom_ptr + 1;  -- increment pointer
                    IF rom_ptr = ROM_SIZE THEN
                        state <= filter0;
                    ELSE
                        state <= config0;
                    END IF;
						
               WHEN filter0 =>
                    if enhance = '1' then
                        z_left <= y_left(0) + x_left(0); -- add output of filter
                        z_right <= y_right(0) + x_right(0); -- to the input
                    else
                        z_left <= x_left(0)(m - 1) & x_left(0); -- input by itself
                        z_right <= x_right(0)(m - 1) & x_right(0); -- pre-pend MSB
                    end if;

                    if (left_right = '0' and left_right_1 = '1') then -- filter runs at the sampling rate
                        x_left(0) := TO_SFIXED(left_in, m - 1, -n); -- convert input vectors to Qm.n format
                        x_right(0) := TO_SFIXED(right_in, m - 1, -n);
                        
                        -- implement IIR left filter
                        acc_left := x_left(0) * b(0) + x_left(1) * b(1) + x_left(2) * b(2) - y_left(1) * a(1) - y_left(2) * a(2); 
                        
                        -- implement IIR right filter
                        acc_right := x_right(0) * b(0) + x_right(1) * b(1) + x_right(2) * b(2) - y_right(1) * a(1) - y_right(2) * a(2);
                        
                        -- update left input delay line
                        x_left(2) := x_left(1);
                        x_left(1) := x_left(0);

                        -- update right input delay line
                        x_right(2) := x_right(1);
                        x_right(1) := x_right(0);

                        -- update left output delay line
                        y_left(0) := acc_left(m - 1 downto -n);
                        y_left(2) := y_left(1);
                        y_left(1) := y_left(0);

                        -- update right output delay line
                        y_right(0) := acc_right(m - 1 downto -n);
                        y_right(2) := y_right(1);
                        y_right(1) := y_right(0);
                    end if;

                    left_out_int <= to_stdlogicvector(z_left); -- convert from SFIXED to std_logic_vector
                    right_out_int <= to_stdlogicvector(z_right); -- convert from SFIXED to std_logic_vector
                    left_out <= left_out_int(m + n - 1 downto 0); -- assign only m+n bits to output vector
                    right_out <= right_out_int(m + n - 1 downto 0); -- assign only m+n bits to output vector
                    left_right_1 <= left_right;
                    state <= filter0;
            END CASE;
        END IF;
    END PROCESS;
END behavioral;